magic
tech scmos
timestamp 1731946603
<< nwell >>
rect -108 -41 110 80
<< ntransistor >>
rect -96 -185 -94 -135
rect -69 -175 -67 -125
rect -44 -170 -42 -145
rect -16 -160 -14 -110
rect 5 -140 7 -124
rect 28 -140 30 -90
rect 49 -112 51 -99
rect 70 -125 72 -75
rect 92 -84 94 -74
<< ptransistor >>
rect -96 -27 -94 73
rect -69 -27 -67 73
rect -44 -27 -42 73
rect -16 23 -14 73
rect 5 -27 7 73
rect 28 40 30 73
rect 49 -27 51 73
rect 70 48 72 73
rect 92 -27 94 73
<< ndiffusion >>
rect -97 -185 -96 -135
rect -94 -185 -93 -135
rect -70 -175 -69 -125
rect -67 -175 -66 -125
rect -45 -170 -44 -145
rect -42 -170 -41 -145
rect -17 -160 -16 -110
rect -14 -160 -13 -110
rect 4 -140 5 -124
rect 7 -140 8 -124
rect 27 -140 28 -90
rect 30 -140 31 -90
rect 48 -112 49 -99
rect 51 -112 52 -99
rect 69 -125 70 -75
rect 72 -125 73 -75
rect 91 -84 92 -74
rect 94 -84 95 -74
<< pdiffusion >>
rect -97 -27 -96 73
rect -94 -27 -93 73
rect -70 -27 -69 73
rect -67 -27 -66 73
rect -45 -27 -44 73
rect -42 -27 -41 73
rect -17 23 -16 73
rect -14 23 -13 73
rect 4 -27 5 73
rect 7 -27 8 73
rect 27 40 28 73
rect 30 40 31 73
rect 48 -27 49 73
rect 51 -27 52 73
rect 69 48 70 73
rect 72 48 73 73
rect 91 -27 92 73
rect 94 -27 95 73
<< ndcontact >>
rect -101 -185 -97 -135
rect -93 -185 -89 -135
rect -74 -175 -70 -125
rect -66 -175 -62 -125
rect -49 -170 -45 -145
rect -41 -170 -37 -145
rect -21 -160 -17 -110
rect -13 -160 -9 -110
rect 0 -140 4 -124
rect 8 -140 12 -124
rect 23 -140 27 -90
rect 31 -140 35 -90
rect 44 -112 48 -99
rect 52 -112 56 -99
rect 65 -125 69 -75
rect 73 -125 77 -75
rect 87 -84 91 -74
rect 95 -84 99 -74
<< pdcontact >>
rect -101 -27 -97 73
rect -93 -27 -89 73
rect -74 -27 -70 73
rect -66 -27 -62 73
rect -49 -27 -45 73
rect -41 -27 -37 73
rect -21 23 -17 73
rect -13 23 -9 73
rect 0 -27 4 73
rect 8 -27 12 73
rect 23 40 27 73
rect 31 40 35 73
rect 44 -27 48 73
rect 52 -27 56 73
rect 65 48 69 73
rect 73 48 77 73
rect 87 -27 91 73
rect 95 -27 99 73
<< polysilicon >>
rect -96 73 -94 76
rect -69 73 -67 76
rect -44 73 -42 76
rect -16 73 -14 76
rect 5 73 7 76
rect 28 73 30 76
rect 49 73 51 76
rect 70 73 72 76
rect 92 73 94 76
rect -96 -135 -94 -27
rect -69 -125 -67 -27
rect -44 -145 -42 -27
rect -16 -110 -14 23
rect 5 -124 7 -27
rect 28 -90 30 40
rect 49 -99 51 -27
rect 70 -75 72 48
rect 92 -74 94 -27
rect 49 -117 51 -112
rect 92 -87 94 -84
rect 70 -129 72 -125
rect 5 -144 7 -140
rect 28 -144 30 -140
rect -16 -164 -14 -160
rect -44 -174 -42 -170
rect -69 -179 -67 -175
rect -96 -189 -94 -185
<< polycontact >>
rect -102 -131 -96 -125
rect -74 -120 -69 -115
rect -48 -111 -44 -106
rect -21 -102 -16 -97
rect 0 -94 5 -89
rect 22 -86 28 -81
rect 43 -78 49 -73
rect 64 -64 70 -59
rect 87 -50 92 -45
<< metal1 >>
rect -108 86 187 94
rect -108 80 110 86
rect -101 73 -97 80
rect -66 73 -62 80
rect -13 73 -9 80
rect 31 73 35 80
rect 73 73 77 80
rect -89 67 -74 73
rect -37 67 -21 73
rect -21 13 -17 23
rect -21 9 0 13
rect 12 67 23 73
rect 23 30 27 40
rect 23 26 44 30
rect 56 67 65 73
rect 65 39 69 48
rect 65 34 87 39
rect 181 31 187 86
rect -74 -34 -70 -27
rect -49 -34 -45 -27
rect -74 -37 -45 -34
rect -148 -50 87 -45
rect 95 -58 99 -27
rect 139 -19 163 -15
rect 209 -19 229 -15
rect 139 -58 143 -19
rect -148 -64 64 -59
rect 87 -62 143 -58
rect -148 -78 43 -73
rect 87 -74 91 -62
rect -148 -86 22 -81
rect -148 -94 0 -89
rect -148 -102 -21 -97
rect -148 -111 -48 -106
rect -148 -120 -74 -115
rect -148 -131 -102 -125
rect -89 -140 -74 -135
rect -49 -138 -21 -134
rect -49 -145 -45 -138
rect -62 -170 -49 -164
rect 0 -115 23 -110
rect 0 -124 4 -115
rect -9 -140 0 -137
rect 44 -93 65 -88
rect 44 -99 48 -93
rect 35 -112 44 -108
rect -101 -193 -97 -185
rect -41 -193 -37 -170
rect 8 -193 12 -140
rect 52 -193 56 -112
rect 77 -84 87 -80
rect 95 -193 99 -84
rect 127 -99 154 -98
rect 170 -99 175 -48
rect 127 -103 175 -99
rect 127 -193 133 -103
rect -126 -204 133 -193
use inv  inv_0
timestamp 1731617906
transform 1 0 170 0 1 3
box -7 -55 39 29
<< labels >>
rlabel metal1 -10 88 -10 88 1 vdd
rlabel metal1 -143 -48 -143 -48 3 g4
rlabel metal1 220 -18 220 -18 1 c4
rlabel metal1 112 -60 112 -60 1 c4bar
rlabel metal1 -142 -62 -142 -62 1 p4
rlabel metal1 -143 -76 -143 -76 3 g3
rlabel metal1 6 -198 6 -198 1 gnd
rlabel metal1 -142 -128 -142 -128 1 c0
rlabel metal1 -142 -118 -142 -118 1 p1
rlabel metal1 -142 -109 -142 -109 1 g1
rlabel metal1 -142 -100 -142 -100 1 p2
rlabel metal1 -143 -92 -143 -92 3 g2
rlabel metal1 -143 -84 -143 -84 3 p3
<< end >>
