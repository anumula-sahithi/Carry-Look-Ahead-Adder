magic
tech scmos
timestamp 1731946245
<< nwell >>
rect -23 -72 166 53
<< ntransistor >>
rect -10 -258 -8 -218
rect 16 -258 18 -218
rect 40 -220 42 -200
rect 60 -244 62 -204
rect 85 -228 87 -215
rect 110 -244 112 -204
rect 137 -223 139 -213
<< ptransistor >>
rect -10 -35 -8 45
rect 16 -35 18 45
rect 40 -35 42 45
rect 60 -6 62 34
rect 85 -35 87 45
rect 110 8 112 34
rect 137 -35 139 45
<< ndiffusion >>
rect -11 -258 -10 -218
rect -8 -258 -7 -218
rect 15 -258 16 -218
rect 18 -258 19 -218
rect 39 -220 40 -200
rect 42 -220 43 -200
rect 59 -244 60 -204
rect 62 -244 63 -204
rect 84 -228 85 -215
rect 87 -228 88 -215
rect 109 -244 110 -204
rect 112 -244 113 -204
rect 136 -223 137 -213
rect 139 -223 140 -213
<< pdiffusion >>
rect -11 -35 -10 45
rect -8 -35 -7 45
rect 15 -35 16 45
rect 18 -35 19 45
rect 39 -35 40 45
rect 42 -35 43 45
rect 59 -6 60 34
rect 62 -6 63 34
rect 84 -35 85 45
rect 87 -35 88 45
rect 109 8 110 34
rect 112 8 113 34
rect 136 -35 137 45
rect 139 -35 140 45
<< ndcontact >>
rect -15 -258 -11 -218
rect -7 -258 -3 -218
rect 11 -258 15 -218
rect 19 -258 23 -218
rect 35 -220 39 -200
rect 43 -220 47 -200
rect 55 -244 59 -204
rect 63 -244 67 -204
rect 80 -228 84 -215
rect 88 -228 92 -215
rect 105 -244 109 -204
rect 113 -244 117 -204
rect 132 -223 136 -213
rect 140 -223 144 -213
<< pdcontact >>
rect -15 -35 -11 45
rect -7 -35 -3 45
rect 11 -35 15 45
rect 19 -35 23 45
rect 35 -35 39 45
rect 43 -35 47 45
rect 55 -6 59 34
rect 63 -6 67 34
rect 80 -35 84 45
rect 88 -35 92 45
rect 105 8 109 34
rect 113 8 117 34
rect 132 -35 136 45
rect 140 -35 144 45
<< polysilicon >>
rect -10 45 -8 48
rect 16 45 18 48
rect 40 45 42 48
rect 60 34 62 48
rect 85 45 87 48
rect -10 -218 -8 -35
rect 16 -218 18 -35
rect 40 -200 42 -35
rect 60 -204 62 -6
rect 110 34 112 48
rect 137 45 139 48
rect -10 -281 -8 -258
rect 16 -280 18 -258
rect 40 -276 42 -220
rect 85 -215 87 -35
rect 110 -204 112 8
rect 137 -167 139 -35
rect 138 -171 139 -167
rect 60 -274 62 -244
rect 85 -270 87 -228
rect 137 -213 139 -171
rect 110 -276 112 -244
rect 137 -273 139 -223
<< polycontact >>
rect -14 -87 -10 -83
rect 12 -101 16 -97
rect 36 -115 40 -111
rect 56 -128 60 -124
rect 81 -141 85 -137
rect 106 -157 110 -153
rect 134 -171 138 -167
<< metal1 >>
rect -23 58 222 63
rect -15 45 -11 58
rect 19 45 23 58
rect -7 -45 -3 -35
rect 11 -45 15 -35
rect 35 -45 39 -35
rect 63 34 67 58
rect 43 -37 47 -35
rect 55 -37 59 -6
rect 43 -41 59 -37
rect -7 -49 39 -45
rect 55 -42 59 -41
rect 80 -42 84 -35
rect 113 34 117 58
rect 88 -38 92 -35
rect 105 -38 109 8
rect 88 -42 109 -38
rect 55 -46 84 -42
rect 105 -43 109 -42
rect 132 -43 136 -35
rect 105 -47 136 -43
rect 216 16 221 58
rect 140 -40 144 -35
rect 175 -35 208 -31
rect 175 -40 181 -35
rect 140 -44 181 -40
rect -64 -87 -14 -83
rect -64 -101 12 -97
rect -64 -115 36 -111
rect -64 -128 56 -124
rect -64 -141 81 -137
rect -65 -157 106 -153
rect -65 -171 134 -167
rect 26 -192 59 -188
rect -15 -290 -11 -258
rect -7 -268 -3 -258
rect 11 -268 15 -258
rect -7 -271 15 -268
rect 19 -266 23 -258
rect 26 -266 30 -192
rect 43 -200 47 -192
rect 19 -270 30 -266
rect 55 -204 59 -192
rect 35 -290 39 -220
rect 63 -196 109 -191
rect 175 -194 181 -44
rect 63 -204 67 -196
rect 88 -215 92 -196
rect 105 -204 109 -196
rect 80 -290 84 -228
rect 113 -199 181 -194
rect 113 -204 117 -199
rect 140 -213 144 -199
rect 132 -290 136 -223
rect 233 -290 242 -65
rect -32 -296 242 -290
rect -32 -297 149 -296
use inv  inv_0
timestamp 1731617906
transform 1 0 215 0 1 -13
box -7 -55 39 29
<< labels >>
rlabel metal1 35 60 35 60 5 vdd
rlabel metal1 5 -47 5 -47 1 k
rlabel metal1 51 -39 51 -39 1 l
rlabel metal1 97 -40 97 -40 1 m
rlabel metal1 -31 -86 -31 -86 1 c0
rlabel metal1 178 -44 178 -44 7 n
rlabel space 252 -32 252 -32 7 c3
rlabel metal1 3 -99 3 -99 1 p1
rlabel metal1 26 -113 26 -113 1 g1
rlabel metal1 49 -126 49 -126 1 p2
rlabel metal1 73 -139 73 -139 1 g2
rlabel metal1 21 -295 21 -295 1 gnd
rlabel metal1 3 -269 3 -269 1 q
rlabel metal1 21 -264 21 -264 1 p
rlabel metal1 79 -194 79 -194 1 o
rlabel metal1 99 -156 99 -156 1 p3
rlabel metal1 126 -170 126 -170 1 g3
<< end >>
