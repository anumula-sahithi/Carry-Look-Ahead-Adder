magic
tech scmos
timestamp 1731946414
<< nwell >>
rect -13 353 62 412
<< ntransistor >>
rect -1 283 1 303
rect 22 283 24 303
rect 49 295 51 305
<< ptransistor >>
rect -1 365 1 405
rect 22 365 24 405
rect 49 365 51 405
<< ndiffusion >>
rect -2 283 -1 303
rect 1 283 2 303
rect 21 283 22 303
rect 24 283 25 303
rect 48 295 49 305
rect 51 295 52 305
<< pdiffusion >>
rect -2 365 -1 405
rect 1 365 2 405
rect 21 365 22 405
rect 24 365 25 405
rect 48 365 49 405
rect 51 365 52 405
<< ndcontact >>
rect -6 283 -2 303
rect 2 283 6 303
rect 17 283 21 303
rect 25 283 29 303
rect 44 295 48 305
rect 52 295 56 305
<< pdcontact >>
rect -6 365 -2 405
rect 2 365 6 405
rect 17 365 21 405
rect 25 365 29 405
rect 44 365 48 405
rect 52 365 56 405
<< polysilicon >>
rect -1 405 1 408
rect 22 405 24 408
rect 49 405 51 408
rect -1 303 1 365
rect 22 303 24 365
rect 49 305 51 365
rect 49 291 51 295
rect -1 277 1 283
rect 22 277 24 283
<< polycontact >>
rect -5 345 -1 349
rect 17 331 22 336
rect 44 316 49 321
<< metal1 >>
rect 102 423 117 429
rect 102 418 106 423
rect -13 414 106 418
rect -13 412 62 414
rect -6 405 -2 412
rect 25 405 29 412
rect 6 400 17 405
rect 17 350 21 365
rect 44 350 48 365
rect -20 345 -5 349
rect 17 346 48 350
rect 102 378 113 382
rect 102 377 107 378
rect -20 331 17 336
rect 52 335 56 365
rect 81 373 107 377
rect 81 335 84 373
rect 143 371 155 379
rect 52 331 84 335
rect -20 316 44 321
rect 52 313 56 331
rect 44 309 56 313
rect 44 305 48 309
rect 6 300 17 303
rect 29 300 44 303
rect 52 289 56 295
rect 115 289 122 346
rect 52 284 122 289
rect -6 272 -2 283
rect 52 272 56 284
rect -6 267 56 272
use inverterl  inverterl_0
timestamp 1731617906
transform 1 0 116 0 1 400
box -7 -55 39 29
<< labels >>
rlabel metal1 -14 347 -14 347 1 c0
rlabel metal1 22 415 22 415 5 vdd
rlabel metal1 149 374 149 374 7 c1
rlabel metal1 -13 333 -13 333 1 p1
rlabel metal1 61 333 61 333 1 c1bar
rlabel metal1 -12 318 -12 318 1 g1
rlabel metal1 25 269 25 269 1 gnd
<< end >>
