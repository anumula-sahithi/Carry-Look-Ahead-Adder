magic
tech scmos
timestamp 1731941149
<< nwell >>
rect 43 -26 81 9
rect 41 -84 79 -45
<< ntransistor >>
rect 131 7 133 17
rect 115 -38 117 -28
<< ptransistor >>
rect 60 -17 62 3
rect 58 -71 60 -51
<< ndiffusion >>
rect 130 7 131 17
rect 133 7 134 17
rect 114 -38 115 -28
rect 117 -38 118 -28
<< pdiffusion >>
rect 59 -17 60 3
rect 62 -17 63 3
rect 57 -71 58 -51
rect 60 -71 61 -51
<< ndcontact >>
rect 126 7 130 17
rect 134 7 138 17
rect 110 -38 114 -28
rect 118 -39 122 -28
<< pdcontact >>
rect 55 -17 59 3
rect 63 -17 67 3
rect 53 -71 57 -51
rect 61 -71 65 -51
<< polysilicon >>
rect 131 17 133 25
rect 60 3 62 13
rect 131 3 133 7
rect 60 -34 62 -17
rect 115 -28 117 0
rect 58 -51 60 -39
rect 115 -56 117 -38
rect 58 -87 60 -71
<< polycontact >>
rect 127 21 131 25
rect 56 -33 60 -29
rect 60 -44 64 -40
rect 111 -55 115 -51
<< metal1 >>
rect 6 63 36 73
rect -43 22 -28 26
rect 10 25 107 26
rect 10 22 127 25
rect -43 -46 -39 22
rect 55 14 96 17
rect 55 3 59 14
rect 6 -11 28 -5
rect 16 -33 56 -29
rect 63 -33 67 -17
rect 16 -46 21 -33
rect 63 -37 75 -33
rect 71 -40 75 -37
rect 64 -44 75 -40
rect 93 -44 96 14
rect 99 -19 103 22
rect 106 21 127 22
rect 99 -23 114 -19
rect 110 -28 114 -23
rect 118 -44 122 -39
rect 126 -33 130 7
rect 126 -42 131 -33
rect -43 -51 21 -46
rect 82 -47 126 -44
rect 61 -51 86 -47
rect 16 -83 21 -51
rect 104 -55 111 -51
rect 104 -62 108 -55
rect 134 -62 138 7
rect 93 -67 138 -62
rect 53 -83 57 -71
rect 16 -87 57 -83
<< m2contact >>
rect 75 -38 80 -33
rect 126 -47 131 -42
rect 88 -67 93 -62
<< metal2 >>
rect 80 -38 92 -33
rect 88 -62 92 -38
rect 131 -47 146 -42
use inverterl  inverterl_0
timestamp 1731617906
transform 1 0 -21 0 1 44
box -7 -55 39 29
<< labels >>
rlabel metal1 28 67 28 67 1 vdd
rlabel metal1 -34 23 -34 23 1 b
rlabel metal1 14 -9 14 -9 1 gnd
rlabel metal1 102 -45 102 -45 1 s
rlabel metal1 107 -64 107 -64 1 a
rlabel metal1 33 23 33 23 1 b_bar
<< end >>
