magic
tech scmos
timestamp 1731949680
<< metal1 >>
rect 163 157 209 162
rect 175 104 241 109
rect -271 78 0 82
rect -271 -143 -268 78
rect -225 64 0 69
rect -202 49 1 54
rect -202 -109 -197 49
rect 142 17 158 21
rect 176 -58 209 -53
rect 200 -104 236 -100
rect -271 -147 -116 -143
rect 140 -147 141 -137
rect -271 -474 -268 -147
rect -225 -155 -95 -154
rect -225 -159 -117 -155
rect -112 -174 -103 -169
rect 140 -176 141 -152
rect -212 -188 -117 -184
rect -212 -189 -64 -188
rect -239 -199 -86 -198
rect -239 -203 -114 -199
rect -239 -339 -234 -203
rect 88 -273 128 -271
rect 133 -273 140 -271
rect 186 -380 209 -375
rect 198 -426 242 -422
rect -271 -478 -119 -474
rect -271 -942 -268 -478
rect -264 -492 -230 -487
rect -225 -492 -115 -487
rect -264 -932 -260 -492
rect -256 -506 -202 -501
rect -197 -506 -113 -501
rect -256 -923 -253 -506
rect -212 -519 -113 -514
rect -234 -532 -111 -527
rect -205 -548 -121 -544
rect -239 -906 -234 -766
rect -205 -898 -201 -548
rect -192 -562 -121 -558
rect -192 -890 -188 -562
rect 190 -791 209 -785
rect 222 -836 230 -832
rect -175 -867 -154 -862
rect -178 -881 -151 -876
rect -192 -895 -150 -890
rect -205 -903 -155 -898
rect -239 -911 -155 -906
rect -212 -919 -150 -914
rect 142 -916 145 -915
rect 150 -916 163 -915
rect -256 -928 -152 -923
rect -264 -937 -149 -932
rect -271 -948 -147 -942
<< m2contact >>
rect 209 157 214 162
rect -230 64 -225 69
rect 118 17 123 22
rect 209 -58 214 -53
rect -202 -114 -197 -109
rect 136 -152 141 -147
rect -230 -159 -225 -154
rect -117 -174 -112 -169
rect -217 -189 -212 -184
rect 128 -273 133 -268
rect -239 -344 -234 -339
rect 209 -380 214 -375
rect 159 -459 166 -450
rect -230 -492 -225 -487
rect -202 -506 -197 -501
rect -217 -519 -212 -514
rect -239 -532 -234 -527
rect -239 -766 -234 -761
rect 145 -687 150 -681
rect 209 -791 214 -785
rect -217 -919 -212 -914
rect 145 -920 150 -915
<< metal2 >>
rect -230 -154 -225 64
rect -239 -527 -234 -344
rect -230 -487 -225 -159
rect -202 -169 -197 -114
rect 118 -147 123 17
rect 209 -53 214 157
rect 118 -152 136 -147
rect -202 -174 -117 -169
rect -239 -761 -234 -532
rect -217 -514 -212 -189
rect -202 -501 -197 -174
rect 128 -450 133 -273
rect 209 -375 214 -58
rect 128 -459 159 -450
rect 128 -461 133 -459
rect -217 -914 -212 -519
rect 145 -915 150 -687
rect 209 -785 214 -380
use val_c4  val_c4_0
timestamp 1731946603
transform 1 0 -7 0 1 -817
box -148 -204 229 94
use val_c3  val_c3_0
timestamp 1731946245
transform 1 0 -56 0 1 -391
box -65 -297 254 63
use val_c2  val_c2_0
timestamp 1731945987
transform 1 0 -4 0 1 -116
box -113 -197 204 93
use val_c1  val_c1_0
timestamp 1731946414
transform 1 0 20 0 1 -267
box -20 267 155 429
<< labels >>
rlabel metal1 230 107 230 107 1 c1
rlabel metal1 200 160 200 160 5 vdd
rlabel metal1 228 -102 228 -102 1 c2
rlabel metal1 232 -424 232 -423 1 c3
rlabel metal1 224 -835 224 -835 1 c4
rlabel metal1 156 19 156 19 1 gnd
rlabel metal1 -153 67 -153 67 1 p1
rlabel metal1 -200 51 -200 51 1 g1
rlabel metal1 -209 -187 -209 -187 1 p2
rlabel metal1 -269 80 -269 80 3 c0
rlabel metal1 -237 -200 -237 -200 1 g2
rlabel metal1 -204 -546 -204 -546 1 p3
rlabel metal1 -189 -562 -189 -562 1 g3
rlabel metal1 -169 -878 -169 -878 1 p4
rlabel metal1 -160 -865 -160 -865 1 g4
<< end >>
