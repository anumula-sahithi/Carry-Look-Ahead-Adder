magic
tech scmos
timestamp 1731617906
<< nwell >>
rect 0 -17 27 20
<< ntransistor >>
rect 13 -35 15 -25
<< ptransistor >>
rect 13 -7 15 13
<< ndiffusion >>
rect 12 -35 13 -25
rect 15 -35 16 -25
<< pdiffusion >>
rect 12 -7 13 13
rect 15 -7 16 13
<< ndcontact >>
rect 8 -35 12 -25
rect 16 -35 20 -25
<< pdcontact >>
rect 8 -7 12 13
rect 16 -7 20 13
<< polysilicon >>
rect 13 13 15 17
rect 13 -25 15 -7
rect 13 -43 15 -35
<< polycontact >>
rect 9 -22 13 -18
<< metal1 >>
rect 0 19 27 29
rect 8 13 12 19
rect 16 -18 20 -7
rect -7 -22 9 -18
rect 16 -22 39 -18
rect 16 -25 20 -22
rect 8 -45 12 -35
rect 0 -55 27 -45
<< labels >>
rlabel metal1 13 25 13 25 5 vdd
rlabel metal1 20 -48 20 -48 1 gnd
rlabel metal1 2 -20 2 -20 1 b
rlabel metal1 29 -20 29 -20 1 Y
<< end >>
