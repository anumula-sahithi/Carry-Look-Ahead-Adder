magic
tech scmos
timestamp 1732063698
<< error_p >>
rect 1461 -26 1467 -25
<< metal1 >>
rect -117 1398 805 1400
rect 1031 1398 1249 1399
rect -117 1395 1305 1398
rect -758 1366 -224 1371
rect -117 1369 -112 1395
rect 800 1379 1305 1395
rect 800 1378 1249 1379
rect -758 1177 -750 1366
rect -211 1159 -206 1163
rect -435 1116 -430 1158
rect 99 1125 108 1313
rect 800 1287 805 1378
rect 909 1232 1048 1237
rect 377 1207 399 1210
rect 426 1119 466 1125
rect 512 1123 518 1133
rect 512 1118 1011 1123
rect -486 1112 -430 1116
rect -757 1105 -739 1109
rect 397 1108 450 1113
rect 522 1110 964 1113
rect 522 1108 599 1110
rect 897 1108 964 1110
rect -212 1038 -206 1042
rect -212 1036 -209 1038
rect -489 985 -483 1036
rect 929 1028 933 1029
rect 903 1024 933 1028
rect -504 981 -483 985
rect -757 964 -751 975
rect 693 956 698 958
rect 693 951 760 956
rect 872 951 940 956
rect 693 944 698 951
rect 427 939 452 944
rect 106 928 121 934
rect -757 828 -751 838
rect -508 780 -502 848
rect -207 775 -201 779
rect 107 769 115 928
rect 107 764 312 769
rect 933 742 940 951
rect 959 912 964 1108
rect 1001 946 1010 1118
rect 1042 961 1048 1232
rect 1295 1069 1305 1379
rect 1295 1061 1898 1069
rect 1295 1015 1305 1061
rect 1887 1028 1897 1061
rect 2263 963 2289 967
rect 1965 955 1982 960
rect 1001 939 1161 946
rect 959 907 1135 912
rect 1129 855 1135 907
rect 1155 885 1161 939
rect 1155 879 1190 885
rect 1290 879 1327 885
rect 1155 878 1161 879
rect 1129 850 1252 855
rect 1290 853 1329 855
rect 1464 853 1468 867
rect 1290 850 1468 853
rect 2264 811 2299 815
rect 1960 803 1977 808
rect 933 736 1027 742
rect -761 686 -754 694
rect -515 675 -508 705
rect 910 702 1248 706
rect 1289 705 1322 710
rect 1031 701 1248 702
rect -210 658 -205 670
rect -210 654 -198 658
rect 1024 596 1032 597
rect 710 591 774 596
rect 864 591 1033 596
rect 710 584 714 591
rect 1024 567 1032 591
rect -764 546 -757 554
rect -517 545 -511 565
rect 105 559 118 563
rect 480 559 485 563
rect 1023 551 1032 567
rect -764 400 -760 406
rect -518 391 -511 417
rect -213 407 -207 539
rect 1023 506 1031 551
rect 1243 438 1248 701
rect 1471 682 1475 699
rect 1290 677 1475 682
rect 2262 658 2300 662
rect 1961 650 1981 655
rect 1290 530 1325 535
rect 1459 506 1463 526
rect 2268 513 2287 517
rect 1312 503 1463 506
rect 1964 505 1987 510
rect 1290 497 1463 503
rect 1243 433 1284 438
rect -213 403 -194 407
rect -213 286 -207 385
rect 442 334 467 339
rect 942 296 950 297
rect 898 292 951 296
rect -512 281 -295 284
rect -213 282 -189 286
rect -522 279 -295 281
rect -763 267 -756 274
rect -763 119 -754 128
rect -514 -73 -510 137
rect -301 136 -295 279
rect 484 261 493 266
rect 484 247 492 252
rect 942 211 950 292
rect 942 206 1202 211
rect 103 198 128 203
rect -301 131 -244 136
rect -249 48 -244 131
rect 1239 124 1246 407
rect 1277 369 1284 433
rect 2273 373 2313 377
rect 1277 365 1303 369
rect 1930 366 1990 370
rect 1463 280 1468 339
rect 1930 211 1935 366
rect 2082 124 2091 336
rect 1239 117 2301 124
rect 51 109 612 114
rect 794 108 2301 117
rect 794 107 877 108
rect 1246 107 2301 108
rect -249 44 -202 48
rect 1461 -28 1467 -26
rect -514 -78 -199 -73
<< m2contact >>
rect -435 1158 -430 1163
rect -217 1158 -211 1163
rect 512 1133 518 1140
rect 99 1119 108 1125
rect 420 1119 426 1125
rect 450 1108 455 1113
rect 516 1108 522 1113
rect -489 1036 -483 1042
rect -217 1036 -212 1042
rect 933 1024 938 1029
rect -529 948 -522 958
rect 760 951 765 956
rect 867 951 872 956
rect 421 939 427 944
rect -508 773 -502 780
rect -213 773 -207 780
rect 312 764 320 769
rect 1042 955 1048 961
rect 1960 955 1965 960
rect 1190 879 1195 885
rect 1284 879 1290 885
rect 1252 850 1257 855
rect 1285 850 1290 855
rect 1955 803 1960 808
rect 1027 736 1033 742
rect 1284 705 1289 710
rect -515 669 -508 675
rect -210 670 -205 675
rect 774 591 779 596
rect -517 539 -511 545
rect -213 539 -207 545
rect 1023 495 1031 506
rect 1285 677 1290 682
rect 1956 650 1961 655
rect 1285 530 1290 535
rect 1959 505 1964 510
rect 1284 497 1290 503
rect 1239 407 1246 412
rect -518 385 -511 391
rect -213 385 -207 391
rect 437 334 442 339
rect 1202 206 1207 211
rect 1930 206 1935 211
<< pdm12contact >>
rect 859 591 864 596
<< metal2 >>
rect -430 1158 -217 1163
rect 438 1133 512 1140
rect 108 1119 420 1125
rect 455 1108 516 1113
rect -797 1101 -791 1106
rect 105 1090 443 1095
rect -483 1036 -217 1042
rect 938 1024 1020 1029
rect -280 958 -272 1004
rect -522 948 -272 958
rect 765 951 867 956
rect 350 938 421 944
rect 351 814 358 938
rect 127 810 358 814
rect 127 808 357 810
rect -502 773 -213 780
rect 127 712 142 808
rect 320 764 433 769
rect 109 706 142 712
rect -508 670 -210 675
rect -508 669 -464 670
rect 1014 620 1019 1024
rect 1863 959 1960 960
rect 1042 867 1048 955
rect 1841 955 1960 959
rect 1841 954 1938 955
rect 1841 901 1847 954
rect 1506 896 1852 901
rect 1195 879 1284 885
rect 1041 842 1048 867
rect 1257 850 1285 855
rect 1041 813 1047 842
rect 1041 806 1264 813
rect 1033 736 1235 742
rect 1229 682 1235 736
rect 1261 710 1264 806
rect 1846 803 1955 808
rect 1846 732 1853 803
rect 1499 727 1853 732
rect 1261 705 1284 710
rect 1229 677 1285 682
rect 1835 650 1956 655
rect 1835 649 1863 650
rect 1014 613 1263 620
rect 779 591 859 596
rect -511 539 -213 545
rect 1258 535 1263 613
rect 1835 556 1844 649
rect 1502 551 1844 556
rect 1258 530 1285 535
rect 1258 529 1263 530
rect 1031 503 1271 506
rect 1810 505 1959 510
rect 1031 497 1284 503
rect 1031 495 1271 497
rect 1246 407 1299 412
rect -511 385 -213 391
rect 1830 375 1841 505
rect 1504 369 1841 375
rect 113 334 437 339
rect 1207 206 1930 211
rect 111 -25 135 -20
rect 128 -26 135 -25
use ff2  ff2_0
timestamp 1732059066
transform 1 0 1973 0 1 920
box -106 -590 301 111
use sum_block  sum_block_0
timestamp 1731961830
transform 1 0 1309 0 1 856
box -34 -527 197 160
use pg_block  pg_block_0
timestamp 1731945508
transform 1 0 -199 0 1 1038
box -81 -1115 312 345
use carry_block  carry_block_0
timestamp 1731949680
transform 1 0 668 0 1 1128
box -271 -1021 242 162
use ff1  ff1_0
timestamp 1732052795
transform 1 0 -710 0 1 1068
box -112 -976 224 112
<< labels >>
rlabel metal1 390 1209 390 1209 1 C0
rlabel metal1 103 1305 103 1305 1 g1
rlabel metal2 113 1093 113 1093 1 p1
rlabel metal1 110 882 110 882 1 g2
rlabel metal2 134 728 134 728 1 p2
rlabel metal1 33 1398 33 1398 5 vdd
rlabel metal1 225 110 225 110 1 gnd
rlabel metal2 140 335 140 335 1 p3
rlabel metal1 482 561 482 561 1 g3
rlabel metal1 110 560 110 560 1 g3
rlabel metal1 487 249 487 249 1 p4
rlabel metal1 490 263 490 263 1 g4
rlabel metal1 116 201 116 201 1 g4
rlabel metal1 915 1234 915 1234 1 c1
rlabel metal1 906 1026 906 1026 1 c2
rlabel metal1 914 705 914 705 1 c3
rlabel metal1 -207 657 -207 657 1 a2
rlabel metal1 -201 404 -201 404 1 b3
rlabel metal1 -203 283 -203 283 1 a3
rlabel metal1 -205 -76 -205 -76 1 a4
rlabel metal2 129 -23 129 -23 1 p4
rlabel metal2 -219 1160 -219 1160 1 b1
rlabel metal1 -752 1107 -752 1107 1 b_1
rlabel metal2 -220 1041 -220 1041 1 a1
rlabel metal1 -754 971 -754 971 1 a_1
rlabel metal2 -217 778 -217 778 1 b2
rlabel metal1 -752 834 -752 834 1 b_2
rlabel metal1 -757 689 -757 689 1 a_2
rlabel metal1 -760 552 -760 552 1 b_3
rlabel metal1 -761 403 -761 403 1 a_3
rlabel metal1 -217 45 -217 45 1 b4
rlabel metal1 -759 124 -759 124 1 a_4
rlabel metal1 -760 270 -760 270 1 b_4
rlabel metal2 -795 1103 -795 1103 1 clk
rlabel metal1 907 294 907 294 1 c_4
rlabel metal2 1510 729 1510 729 1 s_2
rlabel metal2 1514 898 1514 898 1 s_1
rlabel metal2 1526 553 1526 553 1 s_3
rlabel metal2 1520 371 1520 371 1 s_4
rlabel metal1 1464 302 1464 302 1 p4
rlabel space 1946 973 1946 973 1 clk
rlabel metal1 2275 375 2275 375 1 c4
rlabel metal1 2281 515 2281 515 1 s4
rlabel metal1 2276 660 2276 660 1 s3
rlabel metal1 2284 813 2284 813 1 s2
rlabel metal1 2278 965 2278 965 1 s1
<< end >>
